Bit#(8)font[95][12]={
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},/*" ",0*/
{8'h00,8'h00,8'h04,8'h04,8'h04,8'h04,8'h04,8'h04,8'h00,8'h04,8'h00,8'h00},/*"!",1*/
{8'h00,8'h14,8'h0A,8'h0A,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},/*""",2*/
{8'h00,8'h00,8'h14,8'h14,8'h3F,8'h14,8'h0A,8'h3F,8'h0A,8'h0A,8'h00,8'h00},/*"#",3*/
{8'h00,8'h04,8'h1E,8'h15,8'h05,8'h06,8'h0C,8'h14,8'h15,8'h0F,8'h04,8'h00},/*"$",4*/
{8'h00,8'h00,8'h12,8'h15,8'h0D,8'h0A,8'h14,8'h2C,8'h2A,8'h12,8'h00,8'h00},/*"%",5*/
{8'h00,8'h00,8'h04,8'h0A,8'h0A,8'h1E,8'h15,8'h15,8'h09,8'h36,8'h00,8'h00},/*"&",6*/
{8'h00,8'h02,8'h02,8'h01,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},/*"'",7*/
{8'h00,8'h20,8'h10,8'h08,8'h08,8'h08,8'h08,8'h08,8'h08,8'h10,8'h20,8'h00},/*"(",8*/
{8'h00,8'h02,8'h04,8'h08,8'h08,8'h08,8'h08,8'h08,8'h08,8'h04,8'h02,8'h00},/*")",9*/
{8'h00,8'h00,8'h00,8'h04,8'h15,8'h0E,8'h0E,8'h15,8'h04,8'h00,8'h00,8'h00},/*"*",10*/
{8'h00,8'h00,8'h04,8'h04,8'h04,8'h1F,8'h04,8'h04,8'h04,8'h00,8'h00,8'h00},/*"+",11*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h02,8'h02,8'h01},/*",",12*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h1F,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},/*"-",13*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h02,8'h00,8'h00},/*".",14*/
{8'h00,8'h10,8'h08,8'h08,8'h08,8'h04,8'h04,8'h02,8'h02,8'h02,8'h01,8'h00},/*"/",15*/
{8'h00,8'h00,8'h0E,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0E,8'h00,8'h00},/*"0",16*/
{8'h00,8'h00,8'h04,8'h06,8'h04,8'h04,8'h04,8'h04,8'h04,8'h0E,8'h00,8'h00},/*"1",17*/
{8'h00,8'h00,8'h0E,8'h11,8'h11,8'h08,8'h04,8'h02,8'h01,8'h1F,8'h00,8'h00},/*"2",18*/
{8'h00,8'h00,8'h0E,8'h11,8'h10,8'h0C,8'h10,8'h10,8'h11,8'h0E,8'h00,8'h00},/*"3",19*/
{8'h00,8'h00,8'h08,8'h0C,8'h0A,8'h0A,8'h09,8'h1E,8'h08,8'h18,8'h00,8'h00},/*"4",20*/
{8'h00,8'h00,8'h1F,8'h01,8'h01,8'h0F,8'h10,8'h10,8'h11,8'h0E,8'h00,8'h00},/*"5",21*/
{8'h00,8'h00,8'h0E,8'h09,8'h01,8'h0F,8'h11,8'h11,8'h11,8'h0E,8'h00,8'h00},/*"6",22*/
{8'h00,8'h00,8'h1F,8'h09,8'h08,8'h04,8'h04,8'h04,8'h04,8'h04,8'h00,8'h00},/*"7",23*/
{8'h00,8'h00,8'h0E,8'h11,8'h11,8'h0E,8'h11,8'h11,8'h11,8'h0E,8'h00,8'h00},/*"8",24*/
{8'h00,8'h00,8'h0E,8'h11,8'h11,8'h11,8'h1E,8'h10,8'h12,8'h0E,8'h00,8'h00},/*"9",25*/
{8'h00,8'h00,8'h00,8'h00,8'h04,8'h00,8'h00,8'h00,8'h00,8'h04,8'h00,8'h00},/*":",26*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h04,8'h00,8'h00,8'h00,8'h04,8'h04,8'h00},/*";",27*/
{8'h00,8'h20,8'h10,8'h08,8'h04,8'h02,8'h04,8'h08,8'h10,8'h20,8'h00,8'h00},/*"<",28*/
{8'h00,8'h00,8'h00,8'h00,8'h1F,8'h00,8'h00,8'h1F,8'h00,8'h00,8'h00,8'h00},/*"=",29*/
{8'h00,8'h02,8'h04,8'h08,8'h10,8'h20,8'h10,8'h08,8'h04,8'h02,8'h00,8'h00},/*">",30*/
{8'h00,8'h00,8'h0E,8'h11,8'h11,8'h08,8'h04,8'h04,8'h00,8'h04,8'h00,8'h00},/*"?",31*/
{8'h00,8'h00,8'h0E,8'h11,8'h19,8'h15,8'h15,8'h1D,8'h01,8'h1E,8'h00,8'h00},/*"@",32*/
{8'h00,8'h00,8'h04,8'h04,8'h0C,8'h0A,8'h0A,8'h1E,8'h12,8'h33,8'h00,8'h00},/*"A",33*/
{8'h00,8'h00,8'h0F,8'h12,8'h12,8'h0E,8'h12,8'h12,8'h12,8'h0F,8'h00,8'h00},/*"B",34*/
{8'h00,8'h00,8'h1E,8'h11,8'h01,8'h01,8'h01,8'h01,8'h11,8'h0E,8'h00,8'h00},/*"C",35*/
{8'h00,8'h00,8'h0F,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h0F,8'h00,8'h00},/*"D",36*/
{8'h00,8'h00,8'h1F,8'h12,8'h0A,8'h0E,8'h0A,8'h02,8'h12,8'h1F,8'h00,8'h00},/*"E",37*/
{8'h00,8'h00,8'h1F,8'h12,8'h0A,8'h0E,8'h0A,8'h02,8'h02,8'h07,8'h00,8'h00},/*"F",38*/
{8'h00,8'h00,8'h1C,8'h12,8'h01,8'h01,8'h39,8'h11,8'h12,8'h0C,8'h00,8'h00},/*"G",39*/
{8'h00,8'h00,8'h33,8'h12,8'h12,8'h1E,8'h12,8'h12,8'h12,8'h33,8'h00,8'h00},/*"H",40*/
{8'h00,8'h00,8'h1F,8'h04,8'h04,8'h04,8'h04,8'h04,8'h04,8'h1F,8'h00,8'h00},/*"I",41*/
{8'h00,8'h00,8'h3E,8'h08,8'h08,8'h08,8'h08,8'h08,8'h08,8'h09,8'h07,8'h00},/*"J",42*/
{8'h00,8'h00,8'h37,8'h12,8'h0A,8'h06,8'h0A,8'h0A,8'h12,8'h37,8'h00,8'h00},/*"K",43*/
{8'h00,8'h00,8'h07,8'h02,8'h02,8'h02,8'h02,8'h02,8'h22,8'h3F,8'h00,8'h00},/*"L",44*/
{8'h00,8'h00,8'h1B,8'h1B,8'h1B,8'h1B,8'h15,8'h15,8'h15,8'h15,8'h00,8'h00},/*"M",45*/
{8'h00,8'h00,8'h3B,8'h12,8'h16,8'h16,8'h1A,8'h1A,8'h12,8'h17,8'h00,8'h00},/*"N",46*/
{8'h00,8'h00,8'h0E,8'h11,8'h11,8'h11,8'h11,8'h11,8'h11,8'h0E,8'h00,8'h00},/*"O",47*/
{8'h00,8'h00,8'h0F,8'h12,8'h12,8'h0E,8'h02,8'h02,8'h02,8'h07,8'h00,8'h00},/*"P",48*/
{8'h00,8'h00,8'h0E,8'h11,8'h11,8'h11,8'h11,8'h17,8'h19,8'h0E,8'h18,8'h00},/*"Q",49*/
{8'h00,8'h00,8'h0F,8'h12,8'h12,8'h0E,8'h0A,8'h12,8'h12,8'h37,8'h00,8'h00},/*"R",50*/
{8'h00,8'h00,8'h1E,8'h11,8'h01,8'h06,8'h08,8'h10,8'h11,8'h0F,8'h00,8'h00},/*"S",51*/
{8'h00,8'h00,8'h1F,8'h15,8'h04,8'h04,8'h04,8'h04,8'h04,8'h0E,8'h00,8'h00},/*"T",52*/
{8'h00,8'h00,8'h33,8'h12,8'h12,8'h12,8'h12,8'h12,8'h12,8'h0C,8'h00,8'h00},/*"U",53*/
{8'h00,8'h00,8'h33,8'h12,8'h12,8'h0A,8'h0A,8'h0C,8'h04,8'h04,8'h00,8'h00},/*"V",54*/
{8'h00,8'h00,8'h15,8'h15,8'h15,8'h0E,8'h0A,8'h0A,8'h0A,8'h0A,8'h00,8'h00},/*"W",55*/
{8'h00,8'h00,8'h1B,8'h0A,8'h0A,8'h04,8'h04,8'h0A,8'h0A,8'h1B,8'h00,8'h00},/*"X",56*/
{8'h00,8'h00,8'h1B,8'h0A,8'h0A,8'h04,8'h04,8'h04,8'h04,8'h0E,8'h00,8'h00},/*"Y",57*/
{8'h00,8'h00,8'h1F,8'h09,8'h08,8'h04,8'h04,8'h02,8'h12,8'h1F,8'h00,8'h00},/*"Z",58*/
{8'h00,8'h1C,8'h04,8'h04,8'h04,8'h04,8'h04,8'h04,8'h04,8'h04,8'h1C,8'h00},/*"[",59*/
{8'h00,8'h02,8'h02,8'h02,8'h04,8'h04,8'h08,8'h08,8'h08,8'h10,8'h00,8'h00},/*"\",60*/
{8'h00,8'h0E,8'h08,8'h08,8'h08,8'h08,8'h08,8'h08,8'h08,8'h08,8'h0E,8'h00},/*"]",61*/
{8'h00,8'h04,8'h0A,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},/*"^",62*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h3F},/*"_",63*/
{8'h00,8'h04,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00},/*"`",64*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h0C,8'h12,8'h1C,8'h12,8'h3C,8'h00,8'h00},/*"a",65*/
{8'h00,8'h00,8'h03,8'h02,8'h02,8'h0E,8'h12,8'h12,8'h12,8'h0E,8'h00,8'h00},/*"b",66*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h1C,8'h12,8'h02,8'h02,8'h1C,8'h00,8'h00},/*"c",67*/
{8'h00,8'h00,8'h18,8'h10,8'h10,8'h1C,8'h12,8'h12,8'h12,8'h3C,8'h00,8'h00},/*"d",68*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h0C,8'h12,8'h1E,8'h02,8'h1C,8'h00,8'h00},/*"e",69*/
{8'h00,8'h00,8'h38,8'h04,8'h04,8'h1E,8'h04,8'h04,8'h04,8'h1E,8'h00,8'h00},/*"f",70*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h3C,8'h12,8'h0C,8'h02,8'h1E,8'h22,8'h1C},/*"g",71*/
{8'h00,8'h00,8'h03,8'h02,8'h02,8'h0E,8'h12,8'h12,8'h12,8'h37,8'h00,8'h00},/*"h",72*/
{8'h00,8'h00,8'h04,8'h00,8'h00,8'h06,8'h04,8'h04,8'h04,8'h0E,8'h00,8'h00},/*"i",73*/
{8'h00,8'h00,8'h08,8'h00,8'h00,8'h0C,8'h08,8'h08,8'h08,8'h08,8'h08,8'h07},/*"j",74*/
{8'h00,8'h00,8'h03,8'h02,8'h02,8'h3A,8'h0A,8'h0E,8'h12,8'h37,8'h00,8'h00},/*"k",75*/
{8'h00,8'h00,8'h07,8'h04,8'h04,8'h04,8'h04,8'h04,8'h04,8'h1F,8'h00,8'h00},/*"l",76*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h15,8'h15,8'h15,8'h15,8'h00,8'h00},/*"m",77*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h12,8'h12,8'h12,8'h37,8'h00,8'h00},/*"n",78*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h0C,8'h12,8'h12,8'h12,8'h0C,8'h00,8'h00},/*"o",79*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h0F,8'h12,8'h12,8'h12,8'h0E,8'h02,8'h07},/*"p",80*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h1C,8'h12,8'h12,8'h12,8'h1C,8'h10,8'h38},/*"q",81*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h1B,8'h06,8'h02,8'h02,8'h07,8'h00,8'h00},/*"r",82*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h1E,8'h02,8'h0C,8'h10,8'h1E,8'h00,8'h00},/*"s",83*/
{8'h00,8'h00,8'h00,8'h04,8'h04,8'h0E,8'h04,8'h04,8'h04,8'h18,8'h00,8'h00},/*"t",84*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h1B,8'h12,8'h12,8'h12,8'h3C,8'h00,8'h00},/*"u",85*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h37,8'h12,8'h0A,8'h0C,8'h04,8'h00,8'h00},/*"v",86*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h15,8'h15,8'h0E,8'h0A,8'h0A,8'h00,8'h00},/*"w",87*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h1B,8'h0A,8'h04,8'h0A,8'h1B,8'h00,8'h00},/*"x",88*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h37,8'h12,8'h0A,8'h0C,8'h04,8'h04,8'h03},/*"y",89*/
{8'h00,8'h00,8'h00,8'h00,8'h00,8'h1E,8'h08,8'h04,8'h04,8'h1E,8'h00,8'h00},/*"z",90*/
{8'h00,8'h18,8'h08,8'h08,8'h08,8'h04,8'h08,8'h08,8'h08,8'h08,8'h18,8'h00},/*"{",91*/
{8'h08,8'h08,8'h08,8'h08,8'h08,8'h08,8'h08,8'h08,8'h08,8'h08,8'h08,8'h08},/*"|",92*/
{8'h00,8'h06,8'h04,8'h04,8'h04,8'h08,8'h04,8'h04,8'h04,8'h04,8'h06,8'h00},/*"}",93*/
{8'h02,8'h25,8'h18,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00,8'h00}/*"~",94*/
};